//------------------------------------------------------------------------------
// Company: 		 UIUC ECE Dept.
// Engineer:		 Stephen Kempf
//
// Create Date:    
// Design Name:    ECE 385 Lab 5 Given Code - SLC-3 top-level (Physical RAM)
// Module Name:    SLC3
//
// Comments:
//    Revised 03-22-2007
//    Spring 2007 Distribution
//    Revised 07-26-2013
//    Spring 2015 Distribution
//    Revised 09-22-2015 
//    Revised 06-09-2020
//	  Revised 03-02-2021
//------------------------------------------------------------------------------


module slc3(
	input logic [9:0] SW,
	input logic	Clk, Reset, Run, Continue,
	output logic [9:0] LED,
	input logic [15:0] Data_from_SRAM,
	output logic OE, WE,
	output logic [6:0] HEX0, HEX1, HEX2, HEX3,
	output logic [15:0] ADDR,
	output logic [15:0] Data_to_SRAM
);


// An array of 4-bit wires to connect the hex_drivers efficiently to wherever we want
// For Lab 1, they will direclty be connected to the IR register through an always_comb circuit
// For Lab 2, they will be patched into the MEM2IO module so that Memory-mapped IO can take place
logic [3:0] hex_4 [3:0];
logic [3:0] hex_3, hex_2, hex_1, hex_0;



// Internal connections
logic LD_MAR, LD_MDR, LD_IR, LD_BEN, LD_CC, LD_REG, LD_PC, LD_LED;
logic GatePC, GateMDR, GateALU, GateMARMUX;
logic SR2MUX, ADDR1MUX, MARMUX;
logic BEN, MIO_EN, DRMUX, SR1MUX;
logic [1:0] PCMUX, ADDR2MUX, ALUK;
logic [15:0] MDR_In;
logic [15:0] MAR, MDR, IR;




assign hex_3 = IR[15:12];
assign hex_2 = IR[11:8];
assign hex_1 = IR[7:4];
assign hex_0 = IR[3:0];


HexDriver hex_drivers[3:0] ({hex_3, hex_2, hex_1, hex_0}, {HEX3, HEX2, HEX1, HEX0});
// This works thanks to http://stackoverflow.com/questions/1378159/verilog-can-we-have-an-array-of-custom-modules









// Additional internal connections we add
logic [15:0] DataPath_Out;
logic [15:0] PC;
logic [15:0] PC_MUXOUT, MIO_OUT;













// Connect MAR to ADDR, which is also connected as an input into MEM2IO
//	MEM2IO will determine what gets put onto Data_CPU (which serves as a potential
//	input into MDR)
assign ADDR = MAR; 
assign MIO_EN = OE;












//Week 1 registers (MAR, MDR, PC, IR) we add
reg_16 MAR1 (.Clk(Clk), .Load(LD_MAR), .Reset(Reset), .Din(DataPath_Out), .Dout(MAR));
reg_16 MDR1 (.Clk(Clk), .Load(LD_MDR), .Reset(Reset), .Din(MIO_OUT), .Dout(MDR));
reg_16 IR1 (.Clk(Clk), .Load(LD_IR), .Reset(Reset), .Din(DataPath_Out), .Dout(IR));
reg_16 PC1 (.Clk(Clk), .Load(LD_PC), .Reset(Reset), .Din(PC_MUXOUT), .Dout(PC));

//Week 1 multiplexers (PCMUX), MIO_MUX; NEED TO CHANGE IN3
mux4_1 PC_MUX ( .in1(PC+1), .in2(DataPath_Out), .in3(16'b0), .in4(16'bXXXXXXXXXXXXXXXX), .select(PCMUX), .out(PC_MUXOUT));
mux2_1 MIO_MUX ( .in1(MDR_In), .in2(DataPath_Out), .select(MIO_EN), .out(MIO_OUT));
// Connect everything to the data path (you have to figure out this part)
//datapath d0 (.*);
//Our own version of a datapath; NEED TO CHANGE IN1, IN3, IN4
mux16_1 datapath (.in1(16'b0), .in2(PC), .in3(16'b0), .in4(MDR), .select({GateMARMUX, GatePC, GateALU, GateMDR}), .out(DataPath_Out));
















// Our SRAM and I/O controller (note, this plugs into MDR/MAR)
Mem2IO memory_subsystem(
    .*, .Reset(Reset), .ADDR(ADDR), .Switches(SW),
    .HEX0(hex_4[0][3:0]), .HEX1(hex_4[1][3:0]), .HEX2(hex_4[2][3:0]), .HEX3(hex_4[3][3:0]),
    .Data_from_CPU(MDR), .Data_to_CPU(MDR_In),
    .Data_from_SRAM(Data_from_SRAM), .Data_to_SRAM(Data_to_SRAM)
);


// State machine, you need to fill in the code here as well
ISDU state_controller(
	.*, .Reset(Reset), .Run(Run), .Continue(Continue),
	.Opcode(IR[15:12]), .IR_5(IR[5]), .IR_11(IR[11]),
   .Mem_OE(OE), .Mem_WE(WE)
);

// SRAM WE register
//logic SRAM_WE_In, SRAM_WE;
//// SRAM WE synchronizer
//always_ff @(posedge Clk or posedge Reset_ah)
//begin
//	if (Reset_ah) SRAM_WE <= 1'b1; //resets to 1
//	else 
//		SRAM_WE <= SRAM_WE_In;
//end

	
endmodule
